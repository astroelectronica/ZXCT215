.title KiCad schematic
.include "C:/AE/ZXCT215/CEU4J2X7R2A103K125AE_s.mod"
.include "C:/AE/ZXCT215/ZXCT215.LIB"
R1 /IN- /VIN {RSNS}
XU1 /VREF 0 /VSUPPLY /VIN /IN- /CNV ZXCT215
I1 /IN- 0 DC {ILOAD} 
R2 /CNV /OUT {ROUT}
XU2 /OUT 0 CEU4J2X7R2A103K125AE_s
V1 /VIN 0 DC {VIN} 
V3 /VSUPPLY 0 DC {VSUPPLY} 
V2 /VREF 0 DC {VREF} 
.end
